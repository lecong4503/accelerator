module _g (
    input a, b,
    output g
);

assign g = a & b;

endmodule