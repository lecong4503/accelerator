`timescale 1ns / 1ps

module IF_BRAM #(
    parameter DEPTH = 205,
    parameter WIDTH = 40,
    I_F_BW = 8
)
(
    input clk,
    input rst_n,
    input 
)