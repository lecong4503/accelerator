`timescale 1ns / 1ps

module unified_BRAM #(
    parameter I_F_BW = 8,
    parameter W_BW = 8,
    parameter B_BW = 8,
)