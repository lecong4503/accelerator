module and2 (
    input a, b,
    output y
);

assign y = a & b;

endmodule