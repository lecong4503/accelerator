module or2 (
    input a, b,
    output y
);

assign y = a | b;

endmodule